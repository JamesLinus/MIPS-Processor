----------------------------------------------------------------------------------
-- Create Date:    16:38:07 03/09/2016 
-- Module Name:    AND_1Bit - Behavioral 
----------------------------------------------------------------------------------
----------------------------------------------------------------------------------
-- LIBRARIES / PACKAGES
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
----------------------------------------------------------------------------------
-- ENTITY
----------------------------------------------------------------------------------
ENTITY AND_1Bit IS
	PORT(
		a  : IN  STD_LOGIC;
		b  : IN  STD_LOGIC;
		o  : OUT STD_LOGIC 
	);
END AND_1Bit;
----------------------------------------------------------------------------------
-- ARCHITECTURE
----------------------------------------------------------------------------------
ARCHITECTURE Behavioral OF AND_1Bit IS
BEGIN
	o <= a AND b;
END Behavioral;